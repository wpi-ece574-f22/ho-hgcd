module hgcd(
    input wire[7:0] a,
    input wire[7:0] b,
    input wire ld,
    input wire clk,
    input wire reset,
    output wire[7:0] q,
    output wire rdy);

   // design the RTL of this module ..

endmodule
